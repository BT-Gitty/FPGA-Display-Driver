`timescale 1ns / 1ps

module pxl_clock(

    );
endmodule
