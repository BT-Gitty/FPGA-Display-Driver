`timescale 1ns / 1ps

module framebuffer(

/*Practice RTL Memory
    input iClk,
    input iWE,
    input [18:0] iAddr,
    input [11:0] iData,
    output reg [11:0] oData
    );
    
    localparam addrSpace = 307200; //640x480 = 307200
    
    reg [11:0] memory [addrSpace - 1:0];
    
    always @(posedge iClk) begin
        if (iWE) begin
            memory[iAddr] <= iData;
        end
        else begin
            oData <= memory[iAddr];
        end
    end
*/

);

endmodule