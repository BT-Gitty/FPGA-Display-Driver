`timescale 1ns / 1ps

module clock_480(
    input clk_in,
    output clk_out
    
    
    
    );
endmodule
